library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use WORK.micro_pk.all;

package micro_ram_pk is

  constant RAM_CONTENTS : memContents_t (0 to 2 ** ADDR_WIDTH - 1);
  
end package;
------------------------------------------------------------------------------
package body micro_ram_pk is

  constant RAM_CONTENTS : memContents_t (0 to 2 ** ADDR_WIDTH - 1) := (
       0 => "10110000000001000000000000000000",
       1 => "00000000000000000000001000000000",
       2 => "00000000000000000000001000000001",
       3 => "00000000000000000000001000000111",
       4 => "00000000000000000000000000110000",
     512 => "10011000000100000000000000000001",
     513 => "11110000000000001000000000000000",
     514 => "10000000000000000000000000100000",
     515 => "10110000000011000000000000010010",
     516 => "11011000000000000000000000000000",
     517 => "01000000000000000000100000000010",
     518 => "10110000000010000000000000000000",
     519 => "11010000000000000000000000000000",
     520 => "11111000000000000000000000000000",
     521 => "01001000000000000000100000000010",
     522 => "10110000000011000000000000001010",
     523 => "11000000000000000000000000000000",
      others => (others => '0'));
end package body;
